module register_file (
	input CLOCK_50,
	
)